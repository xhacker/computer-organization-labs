`define ALU_AND    3'b000
`define ALU_OR     3'b001
`define ALU_ADD    3'b010
`define ALU_SUB    3'b110
`define ALU_SLT    3'b111